module Subtract(input [15:0] num1, num2, output [15:0] out);
    assign out = num1 - num2;
endmodule